library verilog;
use verilog.vl_types.all;
entity lab5_tb is
end lab5_tb;
